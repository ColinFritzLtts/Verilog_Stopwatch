`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 06/12/2020 11:56:23 AM
// Design Name: 
// Module Name: rtc_displaydriver
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module rtc_displaydriver(
    input [23:0] i_count,
    output [7:0] o_segout1,
    output [7:0] o_segout2,
    output [7:0] o_segout3,
    output [7:0] o_segout4,
    output [7:0] o_segout5,
    output [7:0] o_segout6
    );
endmodule
